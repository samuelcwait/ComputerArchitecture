module not_gate_4bit(x, o);

input [3:0] x;
output [3:0] o;

assign o = ~x;

endmodule
